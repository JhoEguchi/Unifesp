module HD
#(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=12)
(
	input [(DATA_WIDTH-1):0] data,
	input [(ADDR_WIDTH-1):0] addr,
	input we, clk, clk50,
	output reg[(DATA_WIDTH-1):0] q
);

	// Declare the RAM variable
	reg [DATA_WIDTH-1:0] ram[2**ADDR_WIDTH-1:0];

	initial
	begin
	
	ram[0] = 32'b00000111110000000000000000100000;
	ram[1] = 32'b00000111101111100000000000000000;
	ram[2] = 32'b00111000000000000000000110100000;
	ram[3] = 32'b01010011101111110000000000000000;
	ram[4] = 32'b01010011101101000000000000000001;
	ram[5] = 32'b01001000001111010000000000000001;
	ram[6] = 32'b01001000010111010000000000000001;
	ram[7] = 32'b00000100011000100000000000000101;
	ram[8] = 32'b01010100001000110000000000000000;
	ram[9] = 32'b01010011101000010000000000000001;
	ram[10] = 32'b01001000100111010000000000000001;
	ram[11] = 32'b00000011100000000010000000000000;
	ram[12] = 32'b01001011111111010000000000000000;
	ram[13] = 32'b00110111111000000000000000000000;
	ram[14] = 32'b01001011111111010000000000000000;
	ram[15] = 32'b00110111111000000000000000000000;
	ram[16] = 32'b01001000101111010000000000000000;
	ram[17] = 32'b01011000110000000000000000000000;
	ram[18] = 32'b01010100101001100000000000000000;
	ram[19] = 32'b01010011101001010000000000000000;
	ram[20] = 32'b01001000111111010000000000000001;
	ram[21] = 32'b01001100111000000000000000000000;
	ram[22] = 32'b01010011101001110000000000000001;
	ram[23] = 32'b01001001000111010000000000000001;
	ram[24] = 32'b01001000001111010000000000000000;
	ram[25] = 32'b00100100010010000000100000000000;
	ram[26] = 32'b00000111010000000000000000000001;
	ram[27] = 32'b01000100010110100000000110111110;
	ram[28] = 32'b01001000011111010000000000000010;
	ram[29] = 32'b01001000100111010000000000000001;
	ram[30] = 32'b01010110100001000000000000000000;
	ram[31] = 32'b00000111101111010000000000000011;
	ram[32] = 32'b00111100000000000000000110010011;
	ram[33] = 32'b00000000101000001110000000000000;
	ram[34] = 32'b00001111101111010000000000000011;
	ram[35] = 32'b01010100011001010000000000000000;
	ram[36] = 32'b01010011101000110000000000000010;
	ram[37] = 32'b01001000110111010000000000000010;
	ram[38] = 32'b01010110100001100000000000000000;
	ram[39] = 32'b01011100110000000000000000000000;
	ram[40] = 32'b01001000111111010000000000000001;
	ram[41] = 32'b01001001000111010000000000000001;
	ram[42] = 32'b00000100001010000000000000000001;
	ram[43] = 32'b01010100111000010000000000000000;
	ram[44] = 32'b01010011101001110000000000000001;
	ram[45] = 32'b00111000000000000000000110100111;
	ram[46] = 32'b01100100000000000000000000000000;
	ram[128] = 32'b00000111110000000000000000100000;
	ram[129] = 32'b00000111101111100000000000000000;
	ram[130] = 32'b00111000000000000000000111010011;
	ram[131] = 32'b01001000001111010000000000000011;
	ram[132] = 32'b01011000010000000000000000000000;
	ram[133] = 32'b01010100001000100000000000000000;
	ram[134] = 32'b01010011101000010000000000000011;
	ram[135] = 32'b01001000011111010000000000000011;
	ram[136] = 32'b00101000100000110000000000000010;
	ram[137] = 32'b00000111010000000000000000000001;
	ram[138] = 32'b01000100100110100000000111011111;
	ram[139] = 32'b01001000101111010000000000000011;
	ram[140] = 32'b01010110100001010000000000000000;
	ram[141] = 32'b01011100101000000000000000000000;
	ram[142] = 32'b00111000000000000000001000000100;
	ram[143] = 32'b01001000110111010000000000000000;
	ram[144] = 32'b01001100110000000000000000000000;
	ram[145] = 32'b01010011101001100000000000000000;
	ram[146] = 32'b01001000111111010000000000000001;
	ram[147] = 32'b01001100111000000000000000000001;
	ram[148] = 32'b01010011101001110000000000000001;
	ram[149] = 32'b01001001000111010000000000000100;
	ram[150] = 32'b01001101000000000000000000000001;
	ram[151] = 32'b01010011101010000000000000000100;
	ram[152] = 32'b01001000001111010000000000000100;
	ram[153] = 32'b01001000010111010000000000000011;
	ram[154] = 32'b00100100011000010001000000000000;
	ram[155] = 32'b00000111010000000000000000000001;
	ram[156] = 32'b01000100011110100000001000000100;
	ram[157] = 32'b01001000100111010000000000000010;
	ram[158] = 32'b01001000101111010000000000000000;
	ram[159] = 32'b01001000110111010000000000000001;
	ram[160] = 32'b00000000111001010011000000000000;
	ram[161] = 32'b01010100100001110000000000000000;
	ram[162] = 32'b01010011101001000000000000000010;
	ram[163] = 32'b01001001000111010000000000000010;
	ram[164] = 32'b01010110100010000000000000000000;
	ram[165] = 32'b01011101000000000000000000000000;
	ram[166] = 32'b01001000001111010000000000000000;
	ram[167] = 32'b01001000010111010000000000000001;
	ram[168] = 32'b01010100001000100000000000000000;
	ram[169] = 32'b01010011101000010000000000000000;
	ram[170] = 32'b01001000011111010000000000000001;
	ram[171] = 32'b01001000100111010000000000000010;
	ram[172] = 32'b01010100011001000000000000000000;
	ram[173] = 32'b01010011101000110000000000000001;
	ram[174] = 32'b01001000101111010000000000000100;
	ram[175] = 32'b01001000110111010000000000000100;
	ram[176] = 32'b00000100111001100000000000000001;
	ram[177] = 32'b01010100101001110000000000000000;
	ram[178] = 32'b01010011101001010000000000000100;
	ram[179] = 32'b00111000000000000000000111101000;
	ram[180] = 32'b01100100000000000000000000000000;


	end
	
	always @ (negedge clk)
	begin
		// Write
		if (we)
			ram[addr] <= data;
	end

	always @ (negedge clk50)
	begin
		q <= ram[addr];	
	end

endmodule


//module HD (data, address, we, inclock, outclock, q);
//
//	input[31:0] data;
//	input[15:0] address;
//	input we, inclock, outclock;
//	output[31:0] q;
//
//	lpm_ram_dq HDmem(.data(data), .address(address), .we(we), .inclock(inclock), 
//                .outclock(outclock), .q(q));
//	defparam HDmem.lpm_width = 32;
//	defparam HDmem.lpm_widthad = 16;
//	defparam HDmem.lpm_indata = "REGISTERED";
//	defparam HDmem.lpm_outdata = "REGISTERED";
//	defparam HDmem.lpm_file = "hd.mif";
//	
//endmodule