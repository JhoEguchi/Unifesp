module UC(op, sel, oper, writereg, writemem, rjal, smuxjump, smux2beq, out, jump, smux3, smux3beq, controlPC, ls, selectPC, in, smuxdm, smuxreg, smuxHD, writeIM, HDwe, wreReg, smuxAdDM, signalLCD);

	input[5:0] op;
	output reg[1:0] sel, smux3, smux3beq, controlPC, signalLCD;
	output reg[3:0] oper;
	output reg writereg, writemem, rjal, smuxjump, smux2beq, out, jump, ls, selectPC, in, smuxdm, smuxreg, smuxHD, writeIM, HDwe, wreReg, smuxAdDM;
	
	initial
	begin
	signalLCD = 2'b00;
	end
	
	always@ (op) begin
		case(op)
		6'b000000: begin //add
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b10;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b000001: begin //addi
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'b00;
			smux3 = 2'b10;
   		smux3beq = 2'b01;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b000010: begin //sub
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b10;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0001;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b000011: begin //subi
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'b00;
			smux3 = 2'b10;
   		smux3beq = 2'b01;
			controlPC = 2'b00;
			oper = 4'b0001;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b000100: begin //and
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b10;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0010;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b000101: begin //andi
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'b00;
			smux3 = 2'b10;
   		smux3beq = 2'b01;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b000110: begin //or
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b10;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0011;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b000111: begin //ori
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'b00;
			smux3 = 2'b10;
   		smux3beq = 2'b01;
			controlPC = 2'b00;
			oper = 4'b0011;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b001000: begin //not
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b10;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b1001;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b001001: begin //slt
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b10;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b1000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b001010: begin //slti
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'b00;
			smux3 = 2'b10;
   		smux3beq = 2'b01;
			controlPC = 2'b00;
			oper = 4'b1000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b001011: begin //sl
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b10;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0100;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b001100: begin //sr
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b10;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0101;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b001101: begin //jump
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b1;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b01;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b001110: begin //jumpi
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b1;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b1;
			ls = 1'bx;
			sel = 2'b01;
			smux3 = 2'b10;
   		smux3beq = 2'b00;
			controlPC = 2'b01;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b001111: begin //jal
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b1;
			smuxjump = 1'b1;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b1;
			ls = 1'bx;
			sel = 2'b01;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b01;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b010000: begin //beq
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b1;
			smux2beq = 1'b1;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'b00;
			smux3 = 2'b00;
   		smux3beq = 2'b10;
			controlPC = 2'b01;
			oper = 4'b0110;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b010001: begin //bne
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b1;
			smux2beq = 1'b1;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'b00;
			smux3 = 2'b00;
   		smux3beq = 2'b10;
			controlPC = 2'b01;
			oper = 4'b0111;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b010010: begin //load
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'b1;
			sel = 2'b00;
			smux3 = 2'b00;
   		smux3beq = 2'b01;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b010011: begin //loadi
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'b01;
			smux3 = 2'b01;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b010100: begin //store
			writereg = 1'b0;
			writemem = 1'b1;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b1;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'b0;
			sel = 2'b00;
			smux3 = 2'b00;
   		smux3beq = 2'b01;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b010101: begin //move
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b11;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b010110: begin //in
			writereg = 1'b1;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'b10;
			smux3 = 2'b01;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b1;
			in = 1'b1;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = 2'b00;
		end
		6'b010111: begin //out
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b1;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b1;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b011000: begin //nop
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'b0;
			sel = 2'b00;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b011001: begin //hlt
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b10;
   		smux3beq = 2'b00;
			controlPC = 2'b10;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b011100: begin //CpyHDtoIM
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b1;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b011101: begin //CpyRegtoHD
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b1;
			writeIM = 1'b0;
			HDwe = 1'b1;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b011110: begin //CpyHDtoReg
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b1;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b011111: begin //CpyDMtoHD
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b1;
			wreReg = 1'b0;
			smuxAdDM = 1'b1;
			signalLCD = signalLCD;
		end
		6'b100000: begin //CpyHDtoDM
			writereg = 1'b0;
			writemem = 1'b1;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b1;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b1;
			signalLCD = signalLCD;
		end
		6'b100001: begin //TransferToIM
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b100010: begin //displayLCD
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = 2'b01;
		end
		6'b100011: begin //displayPrograma
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = 2'b11;
		end
		6'b100100: begin // setCS
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		6'b100101: begin //unSetCS
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'bx;
			sel = 2'bxx;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end
		default: 
		begin
			writereg = 1'b0;
			writemem = 1'b0;
			rjal = 1'b0;
			smuxjump = 1'b0;
			smux2beq = 1'b0;
			out = 1'b0;
			jump = 1'b0;
			ls = 1'b0;
			sel = 2'b00;
			smux3 = 2'b00;
   		smux3beq = 2'b00;
			controlPC = 2'b00;
			oper = 4'b0000;
			selectPC = 1'b0;
			in = 1'b0;
			smuxdm = 1'b0;
			smuxreg = 1'b0;
			smuxHD = 1'b0;
			writeIM = 1'b0;
			HDwe = 1'b0;
			wreReg = 1'b0;
			smuxAdDM = 1'b0;
			signalLCD = signalLCD;
		end

		endcase
	end
endmodule
	